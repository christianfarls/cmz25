/escnfs/courses/fa24-cse-30342.01/dropbox/dmikolay/VLSI/muddlib.lef